module add (input logic [63:0] a, input logic [63:0] b, output logic [63:0] c);

assign c = a + b;

endmodule
